module ysyx_22050368_exu(




);